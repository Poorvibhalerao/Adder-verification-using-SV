interface intf(input logic clk,input logic reset);
  
  logic [31:0]a;
  logic [31:0] b;
  logic [31:0]out;
  
endinterface;